module hello1();
initial begin
	$display("Hello World");
end
endmodule
